// Controller module for baud and data